`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/06/2024 03:19:38 PM
// Design Name: 
// Module Name: ascii_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mole_rom_ascii(
 input [4:0] row,  // 6-bit row address (0 to 15)
    output reg [63:0] mole_pattern  // 32-bit pattern for each row
);
    always @(*) begin
        case (row)
            5'd0: mole_pattern = 64'b0000000000000000011111111111111111111111111111100000000000000000;  // Row 1
            5'd1: mole_pattern = 64'b0000000000011111111111111111111111111111111111111111100000000000;
            5'd2: mole_pattern = 64'b0000000000011111111111111111111111111111111111111111100000000000;
            5'd3: mole_pattern = 64'b0000000000011111111111111111111111111111111111111111100000000000;
            5'd4: mole_pattern = 64'b0000001111111111111111111111111111111111111111111111111111000000;
            5'd5: mole_pattern = 64'b0000001111111100000011111111111111111111111110000001111111000000;
            5'd6: mole_pattern = 64'b00000011111100001111000111111111111111111111100001100001111000000;
            5'd7: mole_pattern = 64'b0001111111110001110000111111111111111111111100011111001111111000;
            5'd8: mole_pattern = 64'b0001111111110011110000111111111111111111111100111100001111111000;
            5'd9: mole_pattern = 64'b0001111111110011111100111111111111111111111100111111001111111000; // Row 10
            5'd10: mole_pattern = 64'b1111111111100011110001111111111111111111111000111100011111111111; // Row 11
            5'd11: mole_pattern = 64'b111111111111100110011111111111111111111111111001100111111111111; // Row 12
            5'd12: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Row 13
            5'd13: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Row 14
            5'd14: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Row 15
            5'd15: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd16: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd17: mole_pattern = 64'b1111111111111000000000000000000000000000000000000001111111111111; // Blank Row (Row 16)
            5'd18: mole_pattern = 64'b1111111111001111111111111111111111111111111111111100111111111111; // Blank Row (Row 16)
            5'd19: mole_pattern = 64'b1111111100111111111111111111111111111111111111111111001111111111; // Blank Row (Row 16)
            5'd20: mole_pattern = 64'b1111110011111110011111111100000000000000111111111001110011111111; // Blank Row (Row 16)
            5'd21: mole_pattern = 64'b1111110011100111111001111110000000000001111110011111110011111111; // Blank Row (Row 16)
            5'd22: mole_pattern = 64'b1111110011111110011111111111000000000011111111111111110011111111; // Blank Row (Row 16)
            5'd23: mole_pattern = 64'b1111111100111111111111111111100000000111111111100111001111111111; // Blank Row (Row 16)
            5'd24: mole_pattern = 64'b1111111111001111111111111111111111111111111111111100111111111111; // Blank Row (Row 16)
            5'd25: mole_pattern = 64'b1111111111110000000000000000000000000000000000000011111111111111; // Blank Row (Row 16)
            5'd26: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd27: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd28: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd29: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd30: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            5'd31: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Blank Row (Row 16)
            default: mole_pattern = 64'b1111111111111111111111111111111111111111111111111111111111111111; // Default Blank
        endcase
    end
endmodule
